`timescale 1ns / 1ps

// verilator coverage_off
module Buffer_tb (

);
  localparam DELAY_W = 2;
  localparam DATA_W = 1;
  // Inputs
  reg [(DATA_W)-1:0] in0;
  // Outputs
  wire [(DATA_W)-1:0] out0;
  // Control
  reg [(1)-1:0] running;
  reg [(1)-1:0] clk;
  reg [(1)-1:0] rst;
  // Config
  reg [(DELAY_W)-1:0] amount;

  integer i, j;

  localparam CLOCK_PERIOD = 10;

  initial clk = 0;
  always #(CLOCK_PERIOD/2) clk = ~clk;
  `define ADVANCE @(posedge clk) #(CLOCK_PERIOD/2);

  Buffer #(
    .DELAY_W(DELAY_W),
    .DATA_W(DATA_W)
  ) uut (
    .in0(in0),
    .out0(out0),
    .running(running),
    .clk(clk),
    .rst(rst),
    .amount(amount)
  );

  initial begin
    `ifdef VCD;
    $dumpfile("uut.vcd");
    $dumpvars();
    `endif // VCD;
    in0 = 0;
    running = 0;
    clk = 0;
    rst = 0;
    amount = 0;

    `ADVANCE;

    rst = 1;

    `ADVANCE;

    rst = 0;

    `ADVANCE;

    for(i=0;i<(2**DELAY_W);i=i+1) begin
      rst = 1;
      `ADVANCE;
      rst = 0;
      running = 1;
      amount = i[DELAY_W-1:0];
      in0 = i[0];

      `ADVANCE;
      for(j=0;j<i;j=j+1) begin
        `ADVANCE;
      end

      `ADVANCE

      running = 0;
    end

    `ADVANCE;

    amount = 0;

    `ADVANCE;

    $finish();
  end

endmodule
// verilator coverage_on
