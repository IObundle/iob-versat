`timescale 1ns / 1ps

module mem(
	input	clk,
	input	rst, 

	input [31:0] in1,
	input [31:0] in2,
	output reg [31:0] out
	);



endmodule