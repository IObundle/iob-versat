//data and address widths
`define VERSAT_RDATA_W 32
`define VERSAT_WDATA_W 32
`define VERSAT_ADDR_W  26
