`define nYOLO 0
`define nMULADD 1
`include "xyolodefs.vh"
`define PERIOD_W 5
`define nMUL 0
`define DATAPATH_W 16
`define nALULITE 1
`define nBS 0
`define nALU 0
`define nVO 0
`define nMEM 3
`define nSTAGE 5
`define CONF_MEM_ADDR_W 3
`define nVI 0
`define MEM_ADDR_W 5
