`timescale 1ns / 1ps
`include "xversat.vh"

module xreg #(
         parameter DELAY_W = 32,
         parameter ADDR_W = 1,
         parameter DATA_W = 32
              )
    (
    //control
    input                         clk,
    input                         rst,
    
    input                         run,
    output reg                    done,

    // native interface 
    input [DATA_W/8-1:0]          wstrb,
    input [ADDR_W-1:0]            addr,
    input [DATA_W-1:0]            wdata,
    input                         valid,
    output reg                    ready,
    output [DATA_W-1:0]           rdata,

    //input / output data
    input [DATA_W-1:0]            in0,
    output reg [DATA_W-1:0]       out0,

    input [DELAY_W-1:0]           delay0,

    output [DATA_W-1:0]           currentValue
    );

reg [DELAY_W-1:0] delay;
reg running;

assign rdata = (ready ? out0 : 0);
assign currentValue = out0;

always @(posedge clk,posedge rst)
begin
   if(rst) begin
      out0 <= 0;
      delay <= 0;
      ready <= 0;
      done <= 0;
      running <= 0;
   end else begin
      ready <= valid;

      if(valid & |wstrb) begin
         out0 <= wdata;
      end

      if(run) begin
         delay <= delay0;
         running <= 1;
      end 

      if(running) begin
         if(|delay) begin
            delay <= delay - 1;
         end

         if(!done && delay == 0) begin
            out0 <= in0;
            done <= 1;
         end
      end
   end
end

endmodule