
// Versat does not instantiate a testbench unit
